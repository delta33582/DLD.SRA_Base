library verilog;
use verilog.vl_types.all;
entity TEST_COMP_vlg_vec_tst is
end TEST_COMP_vlg_vec_tst;
